// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

module core_ibex_fcov_bind;
  bind ibex_core core_ibex_fcov_bind u_fcov_bind (
    .*
  );
endmodule
